--*****************************************************************************
--***************************  VHDL Source Code  ******************************
--*********  Copyright 2009, Rochester Institute of Technology  ***************
--*****************************************************************************
--
--  DESIGNER NAME:  Bruce Link
--
--       LAB NAME:  cache demo - NIOS based
--
--      FILE NAME:  cache_demo.vhd
--
-------------------------------------------------------------------------------
--
--  DESCRIPTION
--
--    This design is designed to work with the Altera DE1-SoC development board. 
--
--
--  REVISION HISTORY
--
--  _______________________________________________________________________
-- |  DATE    | USER | Ver |  Description                                  |
-- |==========+======+=====+================================================
-- |          |      |     |
-- | 03/01/09 | BAL  | 1.0 | Created
-- |          |      |     |
--
--*****************************************************************************
--*****************************************************************************

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY cache_demo IS
    PORT (
    CLOCK2_50 : IN STD_LOGIC;
    KEY       : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    SW        : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    --
    LEDR    : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) 
        );
END ENTITY cache_demo;

ARCHITECTURE structure OF cache_demo IS

  -----------------------------------------------------------------------------
  -- define components
  -----------------------------------------------------------------------------
  COMPONENT niosSystem IS PORT (
    reset_reset_n         : IN  std_logic;
    clk_clk             : IN  std_logic;
    switches_export : IN  std_logic_vector(7 DOWNTO 0);
    --
    leds_export     : OUT std_logic_vector(7 DOWNTO 0)
  );
  END COMPONENT;

  -----------------------------------------------------------------------------
  -- define custom data types, constants, etc
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  -- define internal signals
  -----------------------------------------------------------------------------

    
BEGIN

    -- Instantiate the Nios II system entity generated by the Qsys Builder
    NiosII : niosSystem PORT MAP (
      clk_clk         => CLOCK2_50,
      reset_reset_n   => KEY(0),
      switches_export => SW,
      --
      leds_export     => LEDR
    );


END ARCHITECTURE Structure;
