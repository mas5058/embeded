// nios_system.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        bus_bridge_acknowledge,    //         bus_bridge.acknowledge
		input  wire        bus_bridge_irq,            //                   .irq
		output wire [10:0] bus_bridge_address,        //                   .address
		output wire        bus_bridge_bus_enable,     //                   .bus_enable
		output wire [3:0]  bus_bridge_byte_enable,    //                   .byte_enable
		output wire        bus_bridge_rw,             //                   .rw
		output wire [31:0] bus_bridge_write_data,     //                   .write_data
		input  wire [31:0] bus_bridge_read_data,      //                   .read_data
		input  wire        clk_clk,                   //                clk.clk
		input  wire [7:0]  eight_bit_input_export,    //    eight_bit_input.export
		output wire        iicclockbit_export,        //        iicclockbit.export
		inout  wire        iicdatabit_export,         //         iicdatabit.export
		input  wire        key1_export,               //               key1.export
		input  wire        reset_reset_n,             //              reset.reset_n
		output wire [15:0] sixteen_bit_output_export  // sixteen_bit_output.export
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                                   // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [16:0] nios2_gen2_0_data_master_address;                                    // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                 // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                       // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                      // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                  // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                            // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                         // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [16:0] nios2_gen2_0_instruction_master_address;                             // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;            // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;         // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;             // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;               // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_chipselect;  // mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_chipselect -> to_external_bus_bridge_0:avalon_chipselect
	wire  [31:0] mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_readdata;    // to_external_bus_bridge_0:avalon_readdata -> mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_readdata
	wire         mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_waitrequest; // to_external_bus_bridge_0:avalon_waitrequest -> mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_waitrequest
	wire   [8:0] mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_address;     // mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_address -> to_external_bus_bridge_0:avalon_address
	wire         mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_read;        // mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_read -> to_external_bus_bridge_0:avalon_read
	wire   [3:0] mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_byteenable;  // mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_byteenable -> to_external_bus_bridge_0:avalon_byteenable
	wire         mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_write;       // mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_write -> to_external_bus_bridge_0:avalon_write
	wire  [31:0] mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_writedata;   // mm_interconnect_0:to_external_bus_bridge_0_avalon_slave_writedata -> to_external_bus_bridge_0:avalon_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;               // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;             // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;          // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;          // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                 // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;            // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_leds_s1_chipselect;                                // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                  // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                   // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                                     // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                 // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_key1_s1_chipselect;                                // mm_interconnect_0:key1_s1_chipselect -> key1:chipselect
	wire  [31:0] mm_interconnect_0_key1_s1_readdata;                                  // key1:readdata -> mm_interconnect_0:key1_s1_readdata
	wire   [1:0] mm_interconnect_0_key1_s1_address;                                   // mm_interconnect_0:key1_s1_address -> key1:address
	wire         mm_interconnect_0_key1_s1_write;                                     // mm_interconnect_0:key1_s1_write -> key1:write_n
	wire  [31:0] mm_interconnect_0_key1_s1_writedata;                                 // mm_interconnect_0:key1_s1_writedata -> key1:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                    // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                      // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;                       // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                    // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                         // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                     // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                         // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_iic_data_bit_s1_chipselect;                        // mm_interconnect_0:iic_data_bit_s1_chipselect -> iic_data_bit:chipselect
	wire  [31:0] mm_interconnect_0_iic_data_bit_s1_readdata;                          // iic_data_bit:readdata -> mm_interconnect_0:iic_data_bit_s1_readdata
	wire   [1:0] mm_interconnect_0_iic_data_bit_s1_address;                           // mm_interconnect_0:iic_data_bit_s1_address -> iic_data_bit:address
	wire         mm_interconnect_0_iic_data_bit_s1_write;                             // mm_interconnect_0:iic_data_bit_s1_write -> iic_data_bit:write_n
	wire  [31:0] mm_interconnect_0_iic_data_bit_s1_writedata;                         // mm_interconnect_0:iic_data_bit_s1_writedata -> iic_data_bit:writedata
	wire         mm_interconnect_0_iic_clock_bit_s1_chipselect;                       // mm_interconnect_0:iic_clock_bit_s1_chipselect -> iic_clock_bit:chipselect
	wire  [31:0] mm_interconnect_0_iic_clock_bit_s1_readdata;                         // iic_clock_bit:readdata -> mm_interconnect_0:iic_clock_bit_s1_readdata
	wire   [1:0] mm_interconnect_0_iic_clock_bit_s1_address;                          // mm_interconnect_0:iic_clock_bit_s1_address -> iic_clock_bit:address
	wire         mm_interconnect_0_iic_clock_bit_s1_write;                            // mm_interconnect_0:iic_clock_bit_s1_write -> iic_clock_bit:write_n
	wire  [31:0] mm_interconnect_0_iic_clock_bit_s1_writedata;                        // mm_interconnect_0:iic_clock_bit_s1_writedata -> iic_clock_bit:writedata
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                                 // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                                  // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         irq_mapper_receiver0_irq;                                            // to_external_bus_bridge_0:avalon_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                            // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                      // rst_controller:reset_out -> [iic_clock_bit:reset_n, iic_data_bit:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, key1:reset_n, leds:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sysid_qsys_0:reset_n, to_external_bus_bridge_0:reset]
	wire         rst_controller_reset_out_reset_req;                                  // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                              // nios2_gen2_0:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                                  // rst_controller_001:reset_out -> [mm_interconnect_0:pio_0_reset_reset_bridge_in_reset_reset, pio_0:reset_n]

	nios_system_iic_clock_bit iic_clock_bit (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_iic_clock_bit_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_iic_clock_bit_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_iic_clock_bit_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_iic_clock_bit_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_iic_clock_bit_s1_readdata),   //                    .readdata
		.out_port   (iicclockbit_export)                             // external_connection.export
	);

	nios_system_iic_data_bit iic_data_bit (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_iic_data_bit_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_iic_data_bit_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_iic_data_bit_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_iic_data_bit_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_iic_data_bit_s1_readdata),   //                    .readdata
		.bidir_port (iicdatabit_export)                             // external_connection.export
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	nios_system_key1 key1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_key1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key1_s1_readdata),   //                    .readdata
		.in_port    (key1_export)                           // external_connection.export
	);

	nios_system_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (sixteen_bit_output_export)             // external_connection.export
	);

	nios_system_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	nios_system_pio_0 pio_0 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_pio_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_0_s1_readdata), //                    .readdata
		.in_port  (eight_bit_input_export)               // external_connection.export
	);

	nios_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_system_to_external_bus_bridge_0 to_external_bus_bridge_0 (
		.clk                (clk_clk),                                                             //                clk.clk
		.reset              (rst_controller_reset_out_reset),                                      //              reset.reset
		.avalon_address     (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_address),     //       avalon_slave.address
		.avalon_byteenable  (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_byteenable),  //                   .byteenable
		.avalon_chipselect  (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_chipselect),  //                   .chipselect
		.avalon_read        (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_read),        //                   .read
		.avalon_write       (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_write),       //                   .write
		.avalon_writedata   (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_writedata),   //                   .writedata
		.avalon_readdata    (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_readdata),    //                   .readdata
		.avalon_waitrequest (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_waitrequest), //                   .waitrequest
		.avalon_irq         (irq_mapper_receiver0_irq),                                            //          interrupt.irq
		.acknowledge        (bus_bridge_acknowledge),                                              // external_interface.export
		.irq                (bus_bridge_irq),                                                      //                   .export
		.address            (bus_bridge_address),                                                  //                   .export
		.bus_enable         (bus_bridge_bus_enable),                                               //                   .export
		.byte_enable        (bus_bridge_byte_enable),                                              //                   .export
		.rw                 (bus_bridge_rw),                                                       //                   .export
		.write_data         (bus_bridge_write_data),                                               //                   .export
		.read_data          (bus_bridge_read_data)                                                 //                   .export
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                     (clk_clk),                                                             //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                                      // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.pio_0_reset_reset_bridge_in_reset_reset           (rst_controller_001_reset_out_reset),                                  //        pio_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                  (nios2_gen2_0_data_master_address),                                    //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest              (nios2_gen2_0_data_master_waitrequest),                                //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable               (nios2_gen2_0_data_master_byteenable),                                 //                                         .byteenable
		.nios2_gen2_0_data_master_read                     (nios2_gen2_0_data_master_read),                                       //                                         .read
		.nios2_gen2_0_data_master_readdata                 (nios2_gen2_0_data_master_readdata),                                   //                                         .readdata
		.nios2_gen2_0_data_master_write                    (nios2_gen2_0_data_master_write),                                      //                                         .write
		.nios2_gen2_0_data_master_writedata                (nios2_gen2_0_data_master_writedata),                                  //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess              (nios2_gen2_0_data_master_debugaccess),                                //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address           (nios2_gen2_0_instruction_master_address),                             //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest       (nios2_gen2_0_instruction_master_waitrequest),                         //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read              (nios2_gen2_0_instruction_master_read),                                //                                         .read
		.nios2_gen2_0_instruction_master_readdata          (nios2_gen2_0_instruction_master_readdata),                            //                                         .readdata
		.iic_clock_bit_s1_address                          (mm_interconnect_0_iic_clock_bit_s1_address),                          //                         iic_clock_bit_s1.address
		.iic_clock_bit_s1_write                            (mm_interconnect_0_iic_clock_bit_s1_write),                            //                                         .write
		.iic_clock_bit_s1_readdata                         (mm_interconnect_0_iic_clock_bit_s1_readdata),                         //                                         .readdata
		.iic_clock_bit_s1_writedata                        (mm_interconnect_0_iic_clock_bit_s1_writedata),                        //                                         .writedata
		.iic_clock_bit_s1_chipselect                       (mm_interconnect_0_iic_clock_bit_s1_chipselect),                       //                                         .chipselect
		.iic_data_bit_s1_address                           (mm_interconnect_0_iic_data_bit_s1_address),                           //                          iic_data_bit_s1.address
		.iic_data_bit_s1_write                             (mm_interconnect_0_iic_data_bit_s1_write),                             //                                         .write
		.iic_data_bit_s1_readdata                          (mm_interconnect_0_iic_data_bit_s1_readdata),                          //                                         .readdata
		.iic_data_bit_s1_writedata                         (mm_interconnect_0_iic_data_bit_s1_writedata),                         //                                         .writedata
		.iic_data_bit_s1_chipselect                        (mm_interconnect_0_iic_data_bit_s1_chipselect),                        //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),             //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),               //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),            //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),           //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),         //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),          //                                         .chipselect
		.key1_s1_address                                   (mm_interconnect_0_key1_s1_address),                                   //                                  key1_s1.address
		.key1_s1_write                                     (mm_interconnect_0_key1_s1_write),                                     //                                         .write
		.key1_s1_readdata                                  (mm_interconnect_0_key1_s1_readdata),                                  //                                         .readdata
		.key1_s1_writedata                                 (mm_interconnect_0_key1_s1_writedata),                                 //                                         .writedata
		.key1_s1_chipselect                                (mm_interconnect_0_key1_s1_chipselect),                                //                                         .chipselect
		.leds_s1_address                                   (mm_interconnect_0_leds_s1_address),                                   //                                  leds_s1.address
		.leds_s1_write                                     (mm_interconnect_0_leds_s1_write),                                     //                                         .write
		.leds_s1_readdata                                  (mm_interconnect_0_leds_s1_readdata),                                  //                                         .readdata
		.leds_s1_writedata                                 (mm_interconnect_0_leds_s1_writedata),                                 //                                         .writedata
		.leds_s1_chipselect                                (mm_interconnect_0_leds_s1_chipselect),                                //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),              //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),                //                                         .write
		.nios2_gen2_0_debug_mem_slave_read                 (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),                 //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),             //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),            //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),           //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),          //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),          //                                         .debugaccess
		.onchip_memory2_0_s1_address                       (mm_interconnect_0_onchip_memory2_0_s1_address),                       //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                         (mm_interconnect_0_onchip_memory2_0_s1_write),                         //                                         .write
		.onchip_memory2_0_s1_readdata                      (mm_interconnect_0_onchip_memory2_0_s1_readdata),                      //                                         .readdata
		.onchip_memory2_0_s1_writedata                     (mm_interconnect_0_onchip_memory2_0_s1_writedata),                     //                                         .writedata
		.onchip_memory2_0_s1_byteenable                    (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                    //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                    (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                    //                                         .chipselect
		.onchip_memory2_0_s1_clken                         (mm_interconnect_0_onchip_memory2_0_s1_clken),                         //                                         .clken
		.pio_0_s1_address                                  (mm_interconnect_0_pio_0_s1_address),                                  //                                 pio_0_s1.address
		.pio_0_s1_readdata                                 (mm_interconnect_0_pio_0_s1_readdata),                                 //                                         .readdata
		.sysid_qsys_0_control_slave_address                (mm_interconnect_0_sysid_qsys_0_control_slave_address),                //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata               (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),               //                                         .readdata
		.to_external_bus_bridge_0_avalon_slave_address     (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_address),     //    to_external_bus_bridge_0_avalon_slave.address
		.to_external_bus_bridge_0_avalon_slave_write       (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_write),       //                                         .write
		.to_external_bus_bridge_0_avalon_slave_read        (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_read),        //                                         .read
		.to_external_bus_bridge_0_avalon_slave_readdata    (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_readdata),    //                                         .readdata
		.to_external_bus_bridge_0_avalon_slave_writedata   (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_writedata),   //                                         .writedata
		.to_external_bus_bridge_0_avalon_slave_byteenable  (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_byteenable),  //                                         .byteenable
		.to_external_bus_bridge_0_avalon_slave_waitrequest (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_waitrequest), //                                         .waitrequest
		.to_external_bus_bridge_0_avalon_slave_chipselect  (mm_interconnect_0_to_external_bus_bridge_0_avalon_slave_chipselect)   //                                         .chipselect
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
